module I2c();

endmodule
